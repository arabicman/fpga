module Complex_Multiplier(input,reset clock);



